module color_rom
	(
		input wire clk,
      input wire [ 7: 0 ] addr,
      output reg [ 23: 0 ] data
	);
	
reg [7 : 0] addr_reg; // address buffer
reg [7 : 0] color;

// Buffering address
always @( posedge clk ) begin
	addr_reg <= addr;
	data <= {color, color, color};
end

// ROM data and declaration
always @( * ) begin
	case ( addr_reg )
		8'h00: color = 8'h00;
		8'h01: color = 8'h01;
		8'h02: color = 8'h02;
		8'h03: color = 8'h03;
		8'h04: color = 8'h04;
		8'h05: color = 8'h05;
		8'h06: color = 8'h06;
		8'h07: color = 8'h07;
		8'h08: color = 8'h08;
		8'h09: color = 8'h09;
		8'h0a: color = 8'h0a;
		8'h0b: color = 8'h0b;
		8'h0c: color = 8'h0c;
		8'h0d: color = 8'h0d;
		8'h0e: color = 8'h0e;
		8'h0f: color = 8'h0f;
		8'h10: color = 8'h10;
		8'h11: color = 8'h11;
		8'h12: color = 8'h12;
		8'h13: color = 8'h13;
		8'h14: color = 8'h14;
		8'h15: color = 8'h15;
		8'h16: color = 8'h16;
		8'h17: color = 8'h17;
		8'h18: color = 8'h18;
		8'h19: color = 8'h19;
		8'h1a: color = 8'h1a;
		8'h1b: color = 8'h1b;
		8'h1c: color = 8'h1c;
		8'h1d: color = 8'h1d;
		8'h1e: color = 8'h1e;
		8'h1f: color = 8'h1f;
		8'h20: color = 8'h20;
		8'h21: color = 8'h21;
		8'h22: color = 8'h22;
		8'h23: color = 8'h23;
		8'h24: color = 8'h24;
		8'h25: color = 8'h25;
		8'h26: color = 8'h26;
		8'h27: color = 8'h27;
		8'h28: color = 8'h28;
		8'h29: color = 8'h29;
		8'h2a: color = 8'h2a;
		8'h2b: color = 8'h2b;
		8'h2c: color = 8'h2c;
		8'h2d: color = 8'h2d;
		8'h2e: color = 8'h2e;
		8'h2f: color = 8'h2f;
		8'h30: color = 8'h30;
		8'h31: color = 8'h31;
		8'h32: color = 8'h32;
		8'h33: color = 8'h33;
		8'h34: color = 8'h34;
		8'h35: color = 8'h35;
		8'h36: color = 8'h36;
		8'h37: color = 8'h37;
		8'h38: color = 8'h38;
		8'h39: color = 8'h39;
		8'h3a: color = 8'h3a;
		8'h3b: color = 8'h3b;
		8'h3c: color = 8'h3c;
		8'h3d: color = 8'h3d;
		8'h3e: color = 8'h3e;
		8'h3f: color = 8'h3f;
		8'h40: color = 8'h40;
		8'h41: color = 8'h41;
		8'h42: color = 8'h42;
		8'h43: color = 8'h43;
		8'h44: color = 8'h44;
		8'h45: color = 8'h45;
		8'h46: color = 8'h46;
		8'h47: color = 8'h47;
		8'h48: color = 8'h48;
		8'h49: color = 8'h49;
		8'h4a: color = 8'h4a;
		8'h4b: color = 8'h4b;
		8'h4c: color = 8'h4c;
		8'h4d: color = 8'h4d;
		8'h4e: color = 8'h4e;
		8'h4f: color = 8'h4f;
		8'h50: color = 8'h50;
		8'h51: color = 8'h51;
		8'h52: color = 8'h52;
		8'h53: color = 8'h53;
		8'h54: color = 8'h54;
		8'h55: color = 8'h55;
		8'h56: color = 8'h56;
		8'h57: color = 8'h57;
		8'h58: color = 8'h58;
		8'h59: color = 8'h59;
		8'h5a: color = 8'h5a;
		8'h5b: color = 8'h5b;
		8'h5c: color = 8'h5c;
		8'h5d: color = 8'h5d;
		8'h5e: color = 8'h5e;
		8'h5f: color = 8'h5f;
		8'h60: color = 8'h60;
		8'h61: color = 8'h61;
		8'h62: color = 8'h62;
		8'h63: color = 8'h63;
		8'h64: color = 8'h64;
		8'h65: color = 8'h65;
		8'h66: color = 8'h66;
		8'h67: color = 8'h67;
		8'h68: color = 8'h68;
		8'h69: color = 8'h69;
		8'h6a: color = 8'h6a;
		8'h6b: color = 8'h6b;
		8'h6c: color = 8'h6c;
		8'h6d: color = 8'h6d;
		8'h6e: color = 8'h6e;
		8'h6f: color = 8'h6f;
		8'h70: color = 8'h70;
		8'h71: color = 8'h71;
		8'h72: color = 8'h72;
		8'h73: color = 8'h73;
		8'h74: color = 8'h74;
		8'h75: color = 8'h75;
		8'h76: color = 8'h76;
		8'h77: color = 8'h77;
		8'h78: color = 8'h78;
		8'h79: color = 8'h79;
		8'h7a: color = 8'h7a;
		8'h7b: color = 8'h7b;
		8'h7c: color = 8'h7c;
		8'h7d: color = 8'h7d;
		8'h7e: color = 8'h7e;
		8'h7f: color = 8'h7f;
		8'h80: color = 8'h80;
		8'h81: color = 8'h81;
		8'h82: color = 8'h82;
		8'h83: color = 8'h83;
		8'h84: color = 8'h84;
		8'h85: color = 8'h85;
		8'h86: color = 8'h86;
		8'h87: color = 8'h87;
		8'h88: color = 8'h88;
		8'h89: color = 8'h89;
		8'h8a: color = 8'h8a;
		8'h8b: color = 8'h8b;
		8'h8c: color = 8'h8c;
		8'h8d: color = 8'h8d;
		8'h8e: color = 8'h8e;
		8'h8f: color = 8'h8f;
		8'h90: color = 8'h90;
		8'h91: color = 8'h91;
		8'h92: color = 8'h92;
		8'h93: color = 8'h93;
		8'h94: color = 8'h94;
		8'h95: color = 8'h95;
		8'h96: color = 8'h96;
		8'h97: color = 8'h97;
		8'h98: color = 8'h98;
		8'h99: color = 8'h99;
		8'h9a: color = 8'h9a;
		8'h9b: color = 8'h9b;
		8'h9c: color = 8'h9c;
		8'h9d: color = 8'h9d;
		8'h9e: color = 8'h9e;
		8'h9f: color = 8'h9f;
		8'ha0: color = 8'ha0;
		8'ha1: color = 8'ha1;
		8'ha2: color = 8'ha2;
		8'ha3: color = 8'ha3;
		8'ha4: color = 8'ha4;
		8'ha5: color = 8'ha5;
		8'ha6: color = 8'ha6;
		8'ha7: color = 8'ha7;
		8'ha8: color = 8'ha8;
		8'ha9: color = 8'ha9;
		8'haa: color = 8'haa;
		8'hab: color = 8'hab;
		8'hac: color = 8'hac;
		8'had: color = 8'had;
		8'hae: color = 8'hae;
		8'haf: color = 8'haf;
		8'hb0: color = 8'hb0;
		8'hb1: color = 8'hb1;
		8'hb2: color = 8'hb2;
		8'hb3: color = 8'hb3;
		8'hb4: color = 8'hb4;
		8'hb5: color = 8'hb5;
		8'hb6: color = 8'hb6;
		8'hb7: color = 8'hb7;
		8'hb8: color = 8'hb8;
		8'hb9: color = 8'hb9;
		8'hba: color = 8'hba;
		8'hbb: color = 8'hbb;
		8'hbc: color = 8'hbc;
		8'hbd: color = 8'hbd;
		8'hbe: color = 8'hbe;
		8'hbf: color = 8'hbf;
		8'hc0: color = 8'hc0;
		8'hc1: color = 8'hc1;
		8'hc2: color = 8'hc2;
		8'hc3: color = 8'hc3;
		8'hc4: color = 8'hc4;
		8'hc5: color = 8'hc5;
		8'hc6: color = 8'hc6;
		8'hc7: color = 8'hc7;
		8'hc8: color = 8'hc8;
		8'hc9: color = 8'hc9;
		8'hca: color = 8'hca;
		8'hcb: color = 8'hcb;
		8'hcc: color = 8'hcc;
		8'hcd: color = 8'hcd;
		8'hce: color = 8'hce;
		8'hcf: color = 8'hcf;
		8'hd0: color = 8'hd0;
		8'hd1: color = 8'hd1;
		8'hd2: color = 8'hd2;
		8'hd3: color = 8'hd3;
		8'hd4: color = 8'hd4;
		8'hd5: color = 8'hd5;
		8'hd6: color = 8'hd6;
		8'hd7: color = 8'hd7;
		8'hd8: color = 8'hd8;
		8'hd9: color = 8'hd9;
		8'hda: color = 8'hda;
		8'hdb: color = 8'hdb;
		8'hdc: color = 8'hdc;
		8'hdd: color = 8'hdd;
		8'hde: color = 8'hde;
		8'hdf: color = 8'hdf;
		8'he0: color = 8'he0;
		8'he1: color = 8'he1;
		8'he2: color = 8'he2;
		8'he3: color = 8'he3;
		8'he4: color = 8'he4;
		8'he5: color = 8'he5;
		8'he6: color = 8'he6;
		8'he7: color = 8'he7;
		8'he8: color = 8'he8;
		8'he9: color = 8'he9;
		8'hea: color = 8'hea;
		8'heb: color = 8'heb;
		8'hec: color = 8'hec;
		8'hed: color = 8'hed;
		8'hee: color = 8'hee;
		8'hef: color = 8'hef;
		8'hf0: color = 8'hf0;
		8'hf1: color = 8'hf1;
		8'hf2: color = 8'hf2;
		8'hf3: color = 8'hf3;
		8'hf4: color = 8'hf4;
		8'hf5: color = 8'hf5;
		8'hf6: color = 8'hf6;
		8'hf7: color = 8'hf7;
		8'hf8: color = 8'hf8;
		8'hf9: color = 8'hf9;
		8'hfa: color = 8'hfa;
		8'hfb: color = 8'hfb;
		8'hfc: color = 8'hfc;
		8'hfd: color = 8'hfd;
		8'hfe: color = 8'hfe;
		8'hff: color = 8'hff;
	endcase
end
	
endmodule