// JRG170, VXS182

/**
 * This module is responsible for converting the serial
 * output from the ADC to the parallel input of the filter
 */
module s2p_conversion
	(
		input shiftin,
		input pout
	);
	
	
endmodule